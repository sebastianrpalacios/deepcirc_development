module gate(_0, _1, _2, _3, _990);
input _0, _1, _2, _3;
output _990;
wire _977, _978, _979, _980, _981, _982, _983, _984, _985, _986, _987;
assign _980 = ~_0;
assign _978 = ~_1;
assign _979 = ~_2;
assign _977 = ~_3;
assign _981 = ~(_2 | _3);
assign _983 = ~(_978 | _980);
assign _984 = ~(_977 | _979);
assign _982 = ~_981;
assign _985 = ~(_983 | _984);
assign _987 = ~(_0 | _982);
assign _986 = ~(_981 | _985);
assign _990 = _986 | _987;
endmodule
