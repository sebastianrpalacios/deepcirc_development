module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _15, _16, _17, _18, _19, _20, _21, _5, _6, _7, _8, _9;
assign _18 = ~_0;
assign _16 = ~_2;
assign _17 = ~_3;
assign _5 = ~(_2 | _3);
assign _8 = ~(_16 | _17);
assign _15 = ~_5;
assign _9 = ~(_5 | _18);
assign _6 = ~(_0 | _15);
assign _19 = ~_9;
assign _7 = ~(_1 | _6);
assign _10 = ~(_8 | _19);
assign _21 = ~_7;
assign _20 = ~_10;
assign _12 = ~(_10 | _21);
assign _11 = ~(_7 | _20);
assign _4 = _11 | _12;
endmodule
