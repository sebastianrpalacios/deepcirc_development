module gate(_0, _1, _2, _3, _1163);
input _0, _1, _2, _3;
output _1163;
wire _1151, _1152, _1153, _1154, _1155, _1156, _1157, _1158, _1159, _1160;
assign _1154 = ~_0;
assign _1153 = ~_1;
assign _1152 = ~_2;
assign _1151 = ~_3;
assign _1155 = ~(_1151 | _1153);
assign _1157 = ~(_2 | _1151);
assign _1159 = ~(_1 | _1151);
assign _1156 = ~(_1152 | _1155);
assign _1158 = ~(_1154 | _1157);
assign _1160 = ~(_1158 | _1159);
assign _1163 = _1156 | _1160;
endmodule
