module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _14, _15, _16, _17, _18, _19, _5, _6, _7, _8, _9;
assign _14 = ~_0;
assign _15 = ~_1;
assign _17 = ~_2;
assign _8 = ~(_1 | _3);
assign _5 = ~(_14 | _15);
assign _7 = ~(_0 | _17);
assign _19 = ~_8;
assign _16 = ~_5;
assign _18 = ~_7;
assign _9 = ~(_7 | _8);
assign _6 = ~(_2 | _16);
assign _10 = ~(_18 | _19);
assign _11 = ~(_9 | _10);
assign _4 = _6 | _11;
endmodule
