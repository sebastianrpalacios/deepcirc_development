module gate(_0, _1, _2, _3, _306);
input _0, _1, _2, _3;
output _306;
wire _298, _299, _300, _301, _302, _303, _304, _305;
assign _298 = ~_0;
assign _299 = ~(_1 | _298);
assign _303 = ~(_2 | _298);
assign _300 = ~(_3 | _299);
assign _301 = ~_300;
assign _304 = ~(_300 | _303);
assign _302 = ~(_2 | _301);
assign _305 = ~(_302 | _304);
assign _306 = _305;
endmodule
