module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _14, _15, _16, _17, _18, _19, _20, _21, _5, _6, _7, _8, _9;
assign _14 = ~_0;
assign _16 = ~_1;
assign _19 = ~_2;
assign _17 = ~_3;
assign _5 = ~(_1 | _14);
assign _7 = ~(_0 | _16);
assign _15 = ~_5;
assign _9 = ~(_5 | _19);
assign _18 = ~_7;
assign _6 = ~(_2 | _15);
assign _20 = ~_9;
assign _8 = ~(_17 | _18);
assign _10 = ~(_7 | _20);
assign _11 = ~(_6 | _8);
assign _21 = ~_11;
assign _4 = _10 | _21;
endmodule
