module gold(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output reg _4;
always @* begin
  {_4} = 1'b0;
  case ({_0, _1, _2, _3})
    4'b0000: {_4} = 1'b1;
    4'b0001: {_4} = 1'b0;
    4'b0010: {_4} = 1'b0;
    4'b0011: {_4} = 1'b1;
    4'b0100: {_4} = 1'b0;
    4'b0101: {_4} = 1'b1;
    4'b0110: {_4} = 1'b1;
    4'b0111: {_4} = 1'b0;
    4'b1000: {_4} = 1'b1;
    4'b1001: {_4} = 1'b1;
    4'b1010: {_4} = 1'b1;
    4'b1011: {_4} = 1'b1;
    4'b1100: {_4} = 1'b0;
    4'b1101: {_4} = 1'b1;
    4'b1110: {_4} = 1'b1;
    4'b1111: {_4} = 1'b1;
  endcase
end
endmodule
