module gate(_0, _1, _2, _3, _819);
input _0, _1, _2, _3;
output _819;
wire _803, _804, _805, _806, _807, _808, _809, _810, _811, _812, _813, _814, _815, _816, _817, _818;
assign _806 = ~_0;
assign _805 = ~_1;
assign _807 = ~(_0 | _1);
assign _804 = ~_2;
assign _803 = ~_3;
assign _810 = ~(_805 | _806);
assign _808 = ~_807;
assign _809 = ~(_3 | _804);
assign _811 = ~(_2 | _803);
assign _812 = ~_811;
assign _813 = ~(_810 | _812);
assign _814 = ~(_809 | _813);
assign _815 = ~_814;
assign _816 = ~(_807 | _814);
assign _817 = ~(_808 | _815);
assign _818 = ~(_816 | _817);
assign _819 = _818;
endmodule
