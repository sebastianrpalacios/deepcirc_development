module gate(_0, _1, _2, _3, _555);
input _0, _1, _2, _3;
output _555;
wire _542, _543, _544, _545, _546, _547, _548, _549, _550, _551, _552, _553, _554;
assign _545 = ~_0;
assign _543 = ~_1;
assign _544 = ~_2;
assign _542 = ~_3;
assign _547 = ~(_1 | _545);
assign _546 = ~(_0 | _543);
assign _551 = ~(_3 | _544);
assign _548 = ~(_544 | _547);
assign _552 = ~(_542 | _547);
assign _549 = ~_548;
assign _553 = ~(_551 | _552);
assign _550 = ~(_546 | _549);
assign _554 = ~(_550 | _553);
assign _555 = _554;
endmodule
