module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _19, _20, _21, _22, _5, _6, _7, _8, _9;
assign _14 = ~_0;
assign _16 = ~_0;
assign _15 = ~_1;
assign _18 = ~_1;
assign _19 = ~_2;
assign _17 = ~_3;
assign _5 = ~(_14 | _15);
assign _8 = ~(_18 | _19);
assign _7 = ~(_16 | _17);
assign _6 = ~(_2 | _5);
assign _20 = ~_8;
assign _21 = ~_6;
assign _9 = ~(_3 | _20);
assign _10 = ~(_7 | _9);
assign _22 = ~_10;
assign _11 = ~(_10 | _21);
assign _12 = ~(_6 | _22);
assign _13 = ~(_11 | _12);
assign _4 = _13;
endmodule
