module gate(_0, _1, _2, _3, _1372);
input _0, _1, _2, _3;
output _1372;
wire _1357, _1358, _1359, _1360, _1361, _1362, _1363, _1364, _1365, _1366, _1367, _1368, _1369, _1370, _1371;
assign _1360 = ~_0;
assign _1359 = ~_1;
assign _1358 = ~_2;
assign _1357 = ~_3;
assign _1364 = ~(_2 | _1360);
assign _1361 = ~(_0 | _1358);
assign _1362 = ~_1361;
assign _1367 = ~(_3 | _1361);
assign _1363 = ~(_1357 | _1362);
assign _1365 = ~(_1363 | _1364);
assign _1368 = ~(_1359 | _1363);
assign _1366 = ~(_1 | _1365);
assign _1369 = ~_1368;
assign _1370 = ~(_1367 | _1369);
assign _1371 = ~(_1366 | _1370);
assign _1372 = _1371;
endmodule
