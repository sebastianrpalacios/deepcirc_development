module gate(_0, _1, _2, _3, _367);
input _0, _1, _2, _3;
output _367;
wire _352, _353, _354, _355, _356, _357, _358, _359, _360, _361, _362, _363, _364, _365, _366;
assign _354 = ~_0;
assign _352 = ~_1;
assign _353 = ~_2;
assign _358 = ~(_2 | _354);
assign _363 = ~(_3 | _352);
assign _355 = ~(_3 | _353);
assign _359 = ~_358;
assign _360 = ~(_1 | _358);
assign _364 = ~_363;
assign _356 = ~_355;
assign _361 = ~_360;
assign _365 = ~(_359 | _364);
assign _357 = ~(_0 | _356);
assign _362 = ~(_357 | _361);
assign _366 = ~(_362 | _365);
assign _367 = _366;
endmodule
