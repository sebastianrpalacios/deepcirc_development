module gate(_0, _1, _2, _3, _155);
input _0, _1, _2, _3;
output _155;
wire _142, _143, _144, _145, _146, _147, _148, _149, _150, _151, _152, _153, _154;
assign _145 = ~_0;
assign _143 = ~_1;
assign _144 = ~_2;
assign _142 = ~_3;
assign _146 = ~(_1 | _145);
assign _149 = ~(_2 | _145);
assign _151 = ~(_0 | _143);
assign _147 = ~(_142 | _146);
assign _152 = ~(_144 | _151);
assign _148 = ~_147;
assign _150 = ~(_147 | _149);
assign _153 = ~(_148 | _152);
assign _154 = ~(_150 | _153);
assign _155 = _154;
endmodule
