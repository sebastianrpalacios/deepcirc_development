module gate(_0, _1, _2, _3, _1277);
input _0, _1, _2, _3;
output _1277;
wire _1261, _1262, _1263, _1264, _1265, _1266, _1267, _1268, _1269, _1270, _1271, _1272, _1273, _1274;
assign _1263 = ~_0;
assign _1261 = ~_1;
assign _1262 = ~_2;
assign _1264 = ~(_3 | _1263);
assign _1267 = ~(_3 | _1262);
assign _1265 = ~(_1261 | _1264);
assign _1268 = ~_1267;
assign _1266 = ~_1265;
assign _1269 = ~(_1265 | _1268);
assign _1270 = ~(_2 | _1266);
assign _1271 = ~(_1269 | _1270);
assign _1272 = ~_1271;
assign _1273 = ~(_1263 | _1271);
assign _1274 = ~(_0 | _1272);
assign _1277 = _1273 | _1274;
endmodule
