module gate(_0, _1, _2, _3, _485);
input _0, _1, _2, _3;
output _485;
wire _473, _474, _475, _476, _477, _478, _479, _480, _481, _482, _483, _484;
assign _475 = ~_0;
assign _474 = ~_2;
assign _473 = ~_3;
assign _476 = ~(_1 | _3);
assign _477 = ~(_1 | _475);
assign _479 = ~(_474 | _476);
assign _478 = ~(_473 | _477);
assign _480 = ~_479;
assign _482 = ~(_476 | _478);
assign _481 = ~(_475 | _480);
assign _483 = ~(_2 | _482);
assign _484 = ~(_481 | _483);
assign _485 = _484;
endmodule
