module gate(_0, _1, _2, _3, _1332);
input _0, _1, _2, _3;
output _1332;
wire _1320, _1321, _1322, _1323, _1324, _1325, _1326, _1327, _1328, _1329, _1330, _1331;
assign _1322 = ~_1;
assign _1321 = ~_2;
assign _1320 = ~_3;
assign _1325 = ~(_1 | _3);
assign _1323 = ~(_0 | _1321);
assign _1328 = ~(_1320 | _1322);
assign _1326 = ~_1325;
assign _1324 = ~_1323;
assign _1329 = ~_1328;
assign _1327 = ~(_1324 | _1326);
assign _1330 = ~(_1323 | _1329);
assign _1331 = ~(_1327 | _1330);
assign _1332 = _1331;
endmodule
