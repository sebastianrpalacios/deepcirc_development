module gate(_0, _1, _2, _3, _1061);
input _0, _1, _2, _3;
output _1061;
wire _1046, _1047, _1048, _1049, _1050, _1051, _1052, _1053, _1054, _1055, _1056, _1057, _1058, _1059, _1060;
assign _1049 = ~_0;
assign _1047 = ~_1;
assign _1048 = ~_2;
assign _1053 = ~(_0 | _2);
assign _1046 = ~_3;
assign _1052 = ~(_2 | _1049);
assign _1050 = ~(_1047 | _1049);
assign _1051 = ~(_1047 | _1048);
assign _1054 = ~(_1 | _1048);
assign _1055 = ~(_1051 | _1052);
assign _1056 = ~(_1053 | _1054);
assign _1057 = ~(_1046 | _1055);
assign _1058 = ~(_3 | _1056);
assign _1059 = ~(_1057 | _1058);
assign _1060 = ~(_1050 | _1059);
assign _1061 = _1060;
endmodule
