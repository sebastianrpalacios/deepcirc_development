module gate(_0, _1, _2, _3, _1260);
input _0, _1, _2, _3;
output _1260;
wire _1248, _1249, _1250, _1251, _1252, _1253, _1254, _1255, _1256, _1257, _1258, _1259;
assign _1250 = ~_0;
assign _1248 = ~_1;
assign _1249 = ~_2;
assign _1251 = ~(_0 | _1248);
assign _1252 = ~(_3 | _1248);
assign _1254 = ~(_1249 | _1251);
assign _1253 = ~(_1250 | _1252);
assign _1255 = ~_1254;
assign _1257 = ~(_1251 | _1253);
assign _1256 = ~(_3 | _1255);
assign _1258 = ~(_2 | _1257);
assign _1259 = ~(_1256 | _1258);
assign _1260 = _1259;
endmodule
