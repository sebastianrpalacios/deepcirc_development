module gate(_0, _1, _2, _3, _845);
input _0, _1, _2, _3;
output _845;
wire _829, _830, _831, _832, _833, _834, _835, _836, _837, _838, _839, _840, _841, _842, _843, _844;
assign _831 = ~_0;
assign _830 = ~_1;
assign _832 = ~_2;
assign _829 = ~_3;
assign _836 = ~(_2 | _3);
assign _833 = ~(_829 | _832);
assign _837 = ~_836;
assign _838 = ~(_1 | _836);
assign _834 = ~(_831 | _833);
assign _841 = ~(_830 | _837);
assign _839 = ~_838;
assign _835 = ~_834;
assign _840 = ~(_835 | _839);
assign _842 = ~(_835 | _841);
assign _843 = ~(_838 | _842);
assign _844 = ~(_840 | _843);
assign _845 = _844;
endmodule
