module gate(_0, _1, _2, _3, _1288);
input _0, _1, _2, _3;
output _1288;
wire _1278, _1279, _1280, _1281, _1282, _1283, _1284, _1285;
assign _1280 = ~(_0 | _1);
assign _1278 = ~_2;
assign _1284 = ~(_2 | _3);
assign _1281 = ~_1280;
assign _1279 = ~(_3 | _1278);
assign _1283 = ~(_0 | _1278);
assign _1282 = ~(_1279 | _1281);
assign _1285 = ~(_1283 | _1284);
assign _1288 = _1282 | _1285;
endmodule
