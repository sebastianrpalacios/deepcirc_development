module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _14, _15, _16, _17, _18, _19, _20, _5, _6, _7, _8, _9;
assign _16 = ~_0;
assign _14 = ~_1;
assign _19 = ~_2;
assign _15 = ~_3;
assign _8 = ~(_2 | _16);
assign _5 = ~(_3 | _14);
assign _10 = ~(_0 | _19);
assign _6 = ~(_1 | _15);
assign _18 = ~_8;
assign _20 = ~_10;
assign _7 = ~(_5 | _6);
assign _17 = ~_7;
assign _11 = ~(_7 | _20);
assign _9 = ~(_17 | _18);
assign _4 = _9 | _11;
endmodule
