module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _15, _16, _17, _18, _19, _20, _5, _6, _7, _8, _9;
assign _15 = ~_0;
assign _19 = ~_1;
assign _20 = ~_1;
assign _17 = ~_2;
assign _16 = ~_3;
assign _10 = ~(_0 | _3);
assign _5 = ~(_15 | _16);
assign _18 = ~_5;
assign _6 = ~(_5 | _17);
assign _7 = ~(_2 | _18);
assign _11 = ~(_6 | _10);
assign _8 = ~(_7 | _19);
assign _12 = ~(_11 | _20);
assign _9 = ~(_6 | _8);
assign _4 = _9 | _12;
endmodule
