module gate(_0, _1, _2, _3, _268);
input _0, _1, _2, _3;
output _268;
wire _260, _261, _262, _263, _264, _265, _266, _267;
assign _260 = ~(_1 | _2);
assign _262 = ~(_0 | _2);
assign _261 = ~_260;
assign _263 = ~(_3 | _262);
assign _264 = ~_263;
assign _266 = ~(_261 | _263);
assign _265 = ~(_260 | _264);
assign _267 = ~(_265 | _266);
assign _268 = _267;
endmodule
