module gate(_0, _1, _2, _3, _1356);
input _0, _1, _2, _3;
output _1356;
wire _1346, _1347, _1348, _1349, _1350, _1351, _1352, _1353, _1354, _1355;
assign _1348 = ~(_0 | _1);
assign _1347 = ~_2;
assign _1346 = ~_3;
assign _1349 = ~(_2 | _3);
assign _1352 = ~(_1346 | _1347);
assign _1350 = ~_1349;
assign _1353 = ~_1352;
assign _1351 = ~(_1348 | _1350);
assign _1354 = ~(_0 | _1353);
assign _1355 = ~(_1351 | _1354);
assign _1356 = _1355;
endmodule
