module m0x32AA (input in2, in1, in4, in3, output out);

	wire \$n6_0;
	wire \$n9_0;
	wire \$n8_0;
	wire \$n7_0;

	nor (\$n7_0, in2, in1);
	not (\$n6_0, in4);
	nor (\$n8_0, \$n6_0, \$n7_0);
	nor (\$n9_0, in1, in3);
	nor (out, \$n9_0, \$n8_0);

endmodule
