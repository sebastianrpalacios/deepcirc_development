module m0x0F (input in2, in1, in3, output out);



endmodule
