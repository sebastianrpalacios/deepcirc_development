module gate(_0, _1, _2, _3, _1422);
input _0, _1, _2, _3;
output _1422;
wire _1408, _1409, _1410, _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421;
assign _1411 = ~_0;
assign _1410 = ~_1;
assign _1409 = ~_2;
assign _1408 = ~_3;
assign _1412 = ~(_1409 | _1411);
assign _1414 = ~(_2 | _1408);
assign _1418 = ~(_1 | _1408);
assign _1413 = ~_1412;
assign _1415 = ~(_1410 | _1414);
assign _1419 = ~_1418;
assign _1416 = ~_1415;
assign _1420 = ~(_1413 | _1419);
assign _1417 = ~(_1412 | _1416);
assign _1421 = ~(_1417 | _1420);
assign _1422 = _1421;
endmodule
