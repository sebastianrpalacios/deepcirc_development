module gate(_0, _1, _2, _3, _1087);
input _0, _1, _2, _3;
output _1087;
wire _1073, _1074, _1075, _1076, _1077, _1078, _1079, _1080, _1081, _1082, _1083, _1084;
assign _1076 = ~_0;
assign _1074 = ~_1;
assign _1075 = ~_2;
assign _1073 = ~_3;
assign _1082 = ~(_1074 | _1076);
assign _1078 = ~(_1 | _1075);
assign _1077 = ~(_1073 | _1076);
assign _1083 = ~(_1073 | _1082);
assign _1079 = ~_1078;
assign _1080 = ~(_1075 | _1077);
assign _1081 = ~(_1077 | _1079);
assign _1084 = ~(_1080 | _1083);
assign _1087 = _1081 | _1084;
endmodule
