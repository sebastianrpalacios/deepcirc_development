module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _19, _20, _21, _22, _23, _24, _25, _26, _27, _28, _5, _6, _7, _8, _9;
assign _22 = ~_0;
assign _23 = ~_0;
assign _25 = ~_1;
assign _19 = ~_2;
assign _24 = ~_2;
assign _20 = ~_3;
assign _6 = ~(_2 | _3);
assign _10 = ~(_23 | _24);
assign _5 = ~(_19 | _20);
assign _21 = ~_6;
assign _11 = ~(_10 | _25);
assign _12 = ~(_0 | _5);
assign _7 = ~(_1 | _21);
assign _27 = ~_11;
assign _26 = ~_12;
assign _8 = ~(_5 | _7);
assign _13 = ~(_6 | _26);
assign _9 = ~(_8 | _22);
assign _28 = ~_13;
assign _14 = ~(_11 | _13);
assign _15 = ~(_27 | _28);
assign _16 = ~(_14 | _15);
assign _4 = _9 | _16;
endmodule
