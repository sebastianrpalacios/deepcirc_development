module gate(_0, _1, _2, _3, _514);
input _0, _1, _2, _3;
output _514;
wire _503, _504, _505, _506, _507, _508, _509, _510, _511, _512, _513;
assign _504 = ~_1;
assign _505 = ~_2;
assign _503 = ~_3;
assign _510 = ~(_0 | _3);
assign _509 = ~(_2 | _504);
assign _506 = ~(_1 | _505);
assign _511 = ~(_509 | _510);
assign _507 = ~(_0 | _506);
assign _512 = ~_511;
assign _508 = ~(_503 | _507);
assign _513 = ~(_508 | _512);
assign _514 = _513;
endmodule
