module m0xCC (input in2, in1, in3, output out);


	not (out, in2);

endmodule
