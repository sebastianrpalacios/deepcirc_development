module gate(_0, _1, _2, _3, _645);
input _0, _1, _2, _3;
output _645;
wire _634, _635, _636, _637, _638, _639, _640, _641, _642;
assign _635 = ~_0;
assign _634 = ~_1;
assign _641 = ~(_1 | _3);
assign _637 = ~(_2 | _635);
assign _636 = ~(_3 | _634);
assign _640 = ~(_2 | _634);
assign _638 = ~_637;
assign _642 = ~(_640 | _641);
assign _639 = ~(_636 | _638);
assign _645 = _639 | _642;
endmodule
