module gate(_0, _1, _2, _3, _883);
input _0, _1, _2, _3;
output _883;
wire _870, _871, _872, _873, _874, _875, _876, _877, _878, _879, _880, _881, _882;
assign _872 = ~_0;
assign _870 = ~_1;
assign _871 = ~_2;
assign _875 = ~(_1 | _2);
assign _880 = ~(_0 | _3);
assign _874 = ~(_3 | _872);
assign _873 = ~(_870 | _871);
assign _879 = ~(_872 | _875);
assign _876 = ~(_874 | _875);
assign _881 = ~(_879 | _880);
assign _877 = ~_876;
assign _878 = ~(_873 | _877);
assign _882 = ~(_878 | _881);
assign _883 = _882;
endmodule
