module gate(_0, _1, _2, _3, _725);
input _0, _1, _2, _3;
output _725;
wire _713, _714, _715, _716, _717, _718, _719, _720, _721, _722, _723, _724;
assign _716 = ~_0;
assign _715 = ~_1;
assign _714 = ~_2;
assign _713 = ~_3;
assign _721 = ~(_1 | _3);
assign _718 = ~(_2 | _715);
assign _717 = ~(_713 | _714);
assign _722 = ~_721;
assign _719 = ~(_717 | _718);
assign _723 = ~(_0 | _722);
assign _720 = ~(_716 | _719);
assign _724 = ~(_720 | _723);
assign _725 = _724;
endmodule
