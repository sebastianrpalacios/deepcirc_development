module gate(_0, _1, _2, _3, _869);
input _0, _1, _2, _3;
output _869;
wire _857, _858, _859, _860, _861, _862, _863, _864, _865, _866, _867, _868;
assign _860 = ~_0;
assign _858 = ~_1;
assign _859 = ~_2;
assign _857 = ~_3;
assign _861 = ~(_2 | _3);
assign _862 = ~(_857 | _859);
assign _863 = ~_862;
assign _865 = ~(_0 | _862);
assign _864 = ~(_860 | _863);
assign _866 = ~(_864 | _865);
assign _867 = ~(_858 | _866);
assign _868 = ~(_861 | _867);
assign _869 = _868;
endmodule
