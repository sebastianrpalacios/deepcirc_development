module gate(_0, _1, _2, _3, _117);
input _0, _1, _2, _3;
output _117;
wire _106, _107, _108, _109, _110, _111, _112, _113, _114, _115, _116;
assign _108 = ~_0;
assign _107 = ~_1;
assign _109 = ~(_1 | _2);
assign _106 = ~_3;
assign _113 = ~(_2 | _108);
assign _110 = ~(_106 | _108);
assign _114 = ~(_107 | _113);
assign _111 = ~_110;
assign _115 = ~(_110 | _114);
assign _112 = ~(_109 | _111);
assign _116 = ~(_112 | _115);
assign _117 = _116;
endmodule
