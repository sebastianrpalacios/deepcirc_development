module gate(_0, _1, _2, _3, _1319);
input _0, _1, _2, _3;
output _1319;
wire _1308, _1309, _1310, _1311, _1312, _1313, _1314, _1315, _1316;
assign _1309 = ~_1;
assign _1308 = ~_3;
assign _1310 = ~(_1 | _3);
assign _1313 = ~(_1308 | _1309);
assign _1311 = ~_1310;
assign _1314 = ~(_0 | _1310);
assign _1312 = ~(_2 | _1311);
assign _1315 = ~_1314;
assign _1316 = ~(_1313 | _1315);
assign _1319 = _1312 | _1316;
endmodule
