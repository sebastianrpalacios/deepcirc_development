module gate(_0, _1, _2, _3, _581);
input _0, _1, _2, _3;
output _581;
wire _568, _569, _570, _571, _572, _573, _574, _575, _576, _577, _578, _579, _580;
assign _571 = ~_0;
assign _569 = ~_1;
assign _570 = ~_2;
assign _568 = ~_3;
assign _574 = ~(_0 | _3);
assign _572 = ~(_568 | _571);
assign _575 = ~(_2 | _574);
assign _573 = ~(_570 | _572);
assign _576 = ~_575;
assign _578 = ~(_569 | _575);
assign _577 = ~(_1 | _576);
assign _579 = ~(_577 | _578);
assign _580 = ~(_573 | _579);
assign _581 = _580;
endmodule
