module gate(_0, _1, _2, _3, _423);
input _0, _1, _2, _3;
output _423;
wire _411, _412, _413, _414, _415, _416, _417, _418, _419, _420, _421, _422;
assign _414 = ~_0;
assign _412 = ~_1;
assign _413 = ~_2;
assign _411 = ~_3;
assign _416 = ~(_3 | _414);
assign _415 = ~(_411 | _412);
assign _417 = ~(_0 | _415);
assign _419 = ~(_415 | _416);
assign _418 = ~_417;
assign _420 = ~(_413 | _419);
assign _421 = ~(_2 | _418);
assign _422 = ~(_420 | _421);
assign _423 = _422;
endmodule
