module gate(_0, _1, _2, _3, _1307);
input _0, _1, _2, _3;
output _1307;
wire _1300, _1301, _1302, _1303, _1304, _1305, _1306;
assign _1301 = ~_0;
assign _1302 = ~(_1 | _2);
assign _1300 = ~_3;
assign _1305 = ~(_3 | _1302);
assign _1303 = ~(_1 | _1300);
assign _1304 = ~(_1301 | _1303);
assign _1306 = ~(_1304 | _1305);
assign _1307 = _1306;
endmodule
