module gate(_0, _1, _2, _3, _229);
input _0, _1, _2, _3;
output _229;
wire _217, _218, _219, _220, _221, _222, _223, _224, _225, _226, _227, _228;
assign _218 = ~_0;
assign _223 = ~(_1 | _2);
assign _217 = ~_3;
assign _222 = ~(_0 | _3);
assign _219 = ~(_217 | _218);
assign _224 = ~(_222 | _223);
assign _220 = ~(_1 | _219);
assign _225 = ~_224;
assign _221 = ~_220;
assign _227 = ~(_220 | _225);
assign _226 = ~(_221 | _224);
assign _228 = ~(_226 | _227);
assign _229 = _228;
endmodule
