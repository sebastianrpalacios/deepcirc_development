module gate(_0, _1, _2, _3, _259);
input _0, _1, _2, _3;
output _259;
wire _249, _250, _251, _252, _253, _254, _255, _256, _257, _258;
assign _250 = ~_1;
assign _249 = ~_3;
assign _253 = ~(_2 | _250);
assign _251 = ~(_1 | _249);
assign _254 = ~(_0 | _253);
assign _252 = ~_251;
assign _255 = ~_254;
assign _256 = ~(_2 | _252);
assign _257 = ~(_251 | _255);
assign _258 = ~(_256 | _257);
assign _259 = _258;
endmodule
