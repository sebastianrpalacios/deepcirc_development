module gate(_0, _1, _2, _3, _389);
input _0, _1, _2, _3;
output _389;
wire _379, _380, _381, _382, _383, _384, _385, _386, _387, _388;
assign _380 = ~_0;
assign _379 = ~_1;
assign _381 = ~_2;
assign _384 = ~(_3 | _379);
assign _382 = ~(_1 | _381);
assign _385 = ~(_380 | _381);
assign _383 = ~(_0 | _382);
assign _386 = ~_385;
assign _387 = ~(_384 | _386);
assign _388 = ~(_383 | _387);
assign _389 = _388;
endmodule
