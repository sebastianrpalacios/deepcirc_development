module gate(_0, _1, _2, _3, _1395);
input _0, _1, _2, _3;
output _1395;
wire _1384, _1385, _1386, _1387, _1388, _1389, _1390, _1391, _1392;
assign _1387 = ~_0;
assign _1386 = ~_1;
assign _1385 = ~_2;
assign _1384 = ~_3;
assign _1388 = ~(_1386 | _1387);
assign _1390 = ~(_1385 | _1386);
assign _1389 = ~(_2 | _1388);
assign _1391 = ~(_1384 | _1390);
assign _1392 = ~_1391;
assign _1395 = _1389 | _1392;
endmodule
