module gate(_0, _1, _2, _3, _746);
input _0, _1, _2, _3;
output _746;
wire _733, _734, _735, _736, _737, _738, _739, _740, _741, _742, _743;
assign _734 = ~_1;
assign _736 = ~(_1 | _2);
assign _733 = ~_3;
assign _735 = ~(_0 | _734);
assign _740 = ~(_2 | _734);
assign _737 = ~(_735 | _736);
assign _741 = ~(_733 | _740);
assign _738 = ~_737;
assign _742 = ~_741;
assign _739 = ~(_3 | _738);
assign _743 = ~(_737 | _742);
assign _746 = _739 | _743;
endmodule
