module gate(_0, _1, _2, _3, _1072);
input _0, _1, _2, _3;
output _1072;
wire _1062, _1063, _1064, _1065, _1066, _1067, _1068, _1069, _1070, _1071;
assign _1063 = ~_1;
assign _1062 = ~_3;
assign _1066 = ~(_2 | _1063);
assign _1064 = ~(_2 | _1062);
assign _1067 = ~(_0 | _1066);
assign _1065 = ~_1064;
assign _1068 = ~_1067;
assign _1070 = ~(_1064 | _1067);
assign _1069 = ~(_1065 | _1068);
assign _1071 = ~(_1069 | _1070);
assign _1072 = _1071;
endmodule
