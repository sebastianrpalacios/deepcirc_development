module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _19, _20, _21, _5, _6, _7, _8, _9;
assign _18 = ~_0;
assign _16 = ~_1;
assign _10 = ~(_0 | _1);
assign _14 = ~_2;
assign _15 = ~_3;
assign _19 = ~_3;
assign _5 = ~(_2 | _3);
assign _20 = ~_10;
assign _6 = ~(_14 | _15);
assign _11 = ~(_19 | _20);
assign _7 = ~(_5 | _6);
assign _17 = ~_7;
assign _9 = ~(_7 | _18);
assign _8 = ~(_16 | _17);
assign _12 = ~(_8 | _11);
assign _21 = ~_12;
assign _13 = ~(_9 | _21);
assign _4 = _13;
endmodule
