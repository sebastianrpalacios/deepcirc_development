module gate(_0, _1, _2, _3, _659);
input _0, _1, _2, _3;
output _659;
wire _646, _647, _648, _649, _650, _651, _652, _653, _654, _655, _656, _657, _658;
assign _649 = ~_0;
assign _648 = ~_1;
assign _647 = ~_2;
assign _646 = ~_3;
assign _650 = ~(_2 | _649);
assign _651 = ~(_0 | _647);
assign _653 = ~(_1 | _650);
assign _652 = ~(_648 | _651);
assign _655 = ~(_651 | _653);
assign _654 = ~(_650 | _652);
assign _657 = ~(_3 | _655);
assign _656 = ~(_646 | _654);
assign _658 = ~(_656 | _657);
assign _659 = _658;
endmodule
