module gate(_0, _1, _2, _3, _919);
input _0, _1, _2, _3;
output _919;
wire _910, _911, _912, _913, _914, _915, _916, _917, _918;
assign _910 = ~_2;
assign _911 = ~(_1 | _3);
assign _915 = ~(_3 | _910);
assign _912 = ~(_2 | _911);
assign _916 = ~(_0 | _915);
assign _913 = ~_912;
assign _917 = ~(_912 | _916);
assign _914 = ~(_0 | _913);
assign _918 = ~(_914 | _917);
assign _919 = _918;
endmodule
