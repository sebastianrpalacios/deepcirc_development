module gate(_0, _1, _2, _3, _436);
input _0, _1, _2, _3;
output _436;
wire _424, _425, _426, _427, _428, _429, _430, _431, _432, _433, _434, _435;
assign _426 = ~_0;
assign _425 = ~_1;
assign _424 = ~_2;
assign _432 = ~(_2 | _426);
assign _427 = ~(_0 | _424);
assign _430 = ~(_1 | _424);
assign _433 = ~(_425 | _432);
assign _428 = ~(_3 | _427);
assign _429 = ~_428;
assign _431 = ~(_428 | _430);
assign _434 = ~(_429 | _433);
assign _435 = ~(_431 | _434);
assign _436 = _435;
endmodule
