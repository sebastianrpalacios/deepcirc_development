module gate(_0, _1, _2, _3, _1133);
input _0, _1, _2, _3;
output _1133;
wire _1120, _1121, _1122, _1123, _1124, _1125, _1126, _1127, _1128, _1129, _1130;
assign _1122 = ~_1;
assign _1121 = ~_2;
assign _1120 = ~_3;
assign _1123 = ~(_2 | _1122);
assign _1126 = ~(_0 | _1120);
assign _1128 = ~(_1120 | _1121);
assign _1124 = ~_1123;
assign _1127 = ~(_1 | _1126);
assign _1125 = ~(_0 | _1124);
assign _1129 = ~(_1127 | _1128);
assign _1130 = ~_1129;
assign _1133 = _1125 | _1130;
endmodule
