module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _13, _14, _15, _5, _6, _7, _8, _9;
assign _6 = ~(_0 | _1);
assign _13 = ~_2;
assign _15 = ~_2;
assign _9 = ~(_2 | _3);
assign _14 = ~_6;
assign _5 = ~(_3 | _13);
assign _8 = ~(_0 | _15);
assign _7 = ~(_5 | _14);
assign _10 = ~(_8 | _9);
assign _4 = _7 | _10;
endmodule
