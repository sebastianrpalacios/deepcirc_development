module gate(_0, _1, _2, _3, _1150);
input _0, _1, _2, _3;
output _1150;
wire _1134, _1135, _1136, _1137, _1138, _1139, _1140, _1141, _1142, _1143, _1144, _1145, _1146, _1147;
assign _1137 = ~_0;
assign _1136 = ~_1;
assign _1135 = ~_2;
assign _1141 = ~(_1 | _2);
assign _1134 = ~_3;
assign _1138 = ~(_1135 | _1136);
assign _1139 = ~_1138;
assign _1140 = ~(_3 | _1138);
assign _1142 = ~(_1134 | _1139);
assign _1143 = ~(_1141 | _1142);
assign _1144 = ~_1143;
assign _1146 = ~(_0 | _1143);
assign _1145 = ~(_1137 | _1144);
assign _1147 = ~(_1145 | _1146);
assign _1150 = _1140 | _1147;
endmodule
