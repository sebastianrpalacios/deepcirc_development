module gate(_0, _1, _2, _3, _472);
input _0, _1, _2, _3;
output _472;
wire _461, _462, _463, _464, _465, _466, _467, _468, _469, _470, _471;
assign _463 = ~_0;
assign _462 = ~_2;
assign _461 = ~_3;
assign _468 = ~(_1 | _3);
assign _464 = ~(_461 | _462);
assign _467 = ~(_0 | _461);
assign _465 = ~(_1 | _464);
assign _469 = ~(_467 | _468);
assign _466 = ~(_463 | _465);
assign _470 = ~(_2 | _469);
assign _471 = ~(_466 | _470);
assign _472 = _471;
endmodule
