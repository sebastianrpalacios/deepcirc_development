module gate(_0, _1, _2, _3, _1001);
input _0, _1, _2, _3;
output _1001;
wire _1000, _991, _992, _993, _994, _995, _996, _997, _998, _999;
assign _991 = ~_1;
assign _995 = ~(_0 | _2);
assign _992 = ~(_0 | _3);
assign _994 = ~(_3 | _991);
assign _993 = ~_992;
assign _996 = ~(_994 | _995);
assign _997 = ~_996;
assign _998 = ~(_992 | _996);
assign _999 = ~(_993 | _997);
assign _1000 = ~(_998 | _999);
assign _1001 = _1000;
endmodule
