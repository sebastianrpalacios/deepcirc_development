module gate(_0, _1, _2, _3, _1011);
input _0, _1, _2, _3;
output _1011;
wire _1002, _1003, _1004, _1005, _1006, _1007, _1008;
assign _1003 = ~_2;
assign _1002 = ~_3;
assign _1004 = ~(_1 | _1003);
assign _1006 = ~(_1002 | _1003);
assign _1005 = ~(_3 | _1004);
assign _1007 = ~(_1 | _1006);
assign _1008 = ~(_0 | _1007);
assign _1011 = _1005 | _1008;
endmodule
