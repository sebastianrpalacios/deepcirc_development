module gate(_0, _1, _2, _3, _1383);
input _0, _1, _2, _3;
output _1383;
wire _1373, _1374, _1375, _1376, _1377, _1378, _1379, _1380;
assign _1375 = ~_0;
assign _1374 = ~_2;
assign _1373 = ~_3;
assign _1379 = ~(_0 | _1374);
assign _1376 = ~(_1373 | _1374);
assign _1377 = ~(_1 | _1376);
assign _1378 = ~(_1375 | _1376);
assign _1380 = ~(_1378 | _1379);
assign _1383 = _1377 | _1380;
endmodule
