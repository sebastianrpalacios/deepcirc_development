module gate(_0, _1, _2, _3, _976);
input _0, _1, _2, _3;
output _976;
wire _959, _960, _961, _962, _963, _964, _965, _966, _967, _968, _969, _970, _971, _972, _973, _974, _975;
assign _961 = ~_1;
assign _960 = ~_2;
assign _959 = ~_3;
assign _968 = ~(_3 | _961);
assign _971 = ~(_0 | _960);
assign _962 = ~(_0 | _959);
assign _964 = ~(_959 | _961);
assign _965 = ~(_1 | _959);
assign _972 = ~_971;
assign _963 = ~(_1 | _962);
assign _966 = ~_965;
assign _969 = ~(_963 | _964);
assign _967 = ~(_0 | _966);
assign _973 = ~(_969 | _972);
assign _970 = ~(_967 | _968);
assign _974 = ~(_2 | _970);
assign _975 = ~(_973 | _974);
assign _976 = _975;
endmodule
