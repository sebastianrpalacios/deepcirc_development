module gate(_0, _1, _2, _3, _1247);
input _0, _1, _2, _3;
output _1247;
wire _1231, _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243, _1244, _1245, _1246;
assign _1234 = ~_0;
assign _1233 = ~_1;
assign _1232 = ~_2;
assign _1231 = ~_3;
assign _1242 = ~(_2 | _1234);
assign _1235 = ~(_2 | _1233);
assign _1239 = ~(_3 | _1233);
assign _1236 = ~(_1231 | _1234);
assign _1243 = ~_1242;
assign _1237 = ~_1236;
assign _1238 = ~(_1235 | _1237);
assign _1240 = ~(_1238 | _1239);
assign _1241 = ~_1240;
assign _1245 = ~(_1240 | _1243);
assign _1244 = ~(_1232 | _1241);
assign _1246 = ~(_1244 | _1245);
assign _1247 = _1246;
endmodule
