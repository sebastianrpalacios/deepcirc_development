module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _15, _16, _17, _18, _19, _20, _21, _22, _5, _6, _7, _8, _9;
assign _16 = ~_0;
assign _19 = ~_0;
assign _18 = ~_1;
assign _15 = ~_2;
assign _20 = ~_3;
assign _8 = ~(_0 | _3);
assign _7 = ~(_2 | _18);
assign _5 = ~(_1 | _15);
assign _9 = ~(_19 | _20);
assign _17 = ~_5;
assign _10 = ~(_5 | _7);
assign _11 = ~(_8 | _9);
assign _6 = ~(_16 | _17);
assign _21 = ~_10;
assign _22 = ~_11;
assign _12 = ~(_21 | _22);
assign _4 = _6 | _12;
endmodule
