module gate(_0, _1, _2, _3, _948);
input _0, _1, _2, _3;
output _948;
wire _933, _934, _935, _936, _937, _938, _939, _940, _941, _942, _943, _944, _945, _946, _947;
assign _935 = ~_0;
assign _933 = ~_1;
assign _934 = ~_2;
assign _936 = ~(_1 | _3);
assign _941 = ~(_2 | _933);
assign _938 = ~(_0 | _934);
assign _937 = ~_936;
assign _942 = ~_941;
assign _939 = ~_938;
assign _944 = ~(_936 | _938);
assign _943 = ~(_935 | _942);
assign _940 = ~(_937 | _939);
assign _945 = ~_944;
assign _946 = ~(_943 | _945);
assign _947 = ~(_940 | _946);
assign _948 = _947;
endmodule
