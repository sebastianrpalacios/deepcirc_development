module gate(_0, _1, _2, _3, _909);
input _0, _1, _2, _3;
output _909;
wire _898, _899, _900, _901, _902, _903, _904, _905, _906, _907, _908;
assign _899 = ~_0;
assign _898 = ~_2;
assign _900 = ~(_2 | _899);
assign _902 = ~(_0 | _898);
assign _901 = ~_900;
assign _903 = ~(_3 | _902);
assign _904 = ~(_1 | _903);
assign _905 = ~_904;
assign _907 = ~(_901 | _904);
assign _906 = ~(_900 | _905);
assign _908 = ~(_906 | _907);
assign _909 = _908;
endmodule
