module m0xF0 (input in2, in1, in3, output out);


	not (out, in1);

endmodule
