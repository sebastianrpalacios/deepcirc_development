module gate(_0, _1, _2, _3, _787);
input _0, _1, _2, _3;
output _787;
wire _775, _776, _777, _778, _779, _780, _781, _782, _783, _784, _785, _786;
assign _776 = ~_1;
assign _777 = ~_2;
assign _775 = ~_3;
assign _778 = ~(_2 | _3);
assign _781 = ~(_3 | _776);
assign _783 = ~(_775 | _777);
assign _779 = ~(_0 | _778);
assign _784 = ~(_1 | _783);
assign _780 = ~_779;
assign _782 = ~(_779 | _781);
assign _785 = ~(_780 | _784);
assign _786 = ~(_782 | _785);
assign _787 = _786;
endmodule
