module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _5, _6, _7, _8, _9;
assign _15 = ~_0;
assign _5 = ~(_0 | _1);
assign _13 = ~_2;
assign _16 = ~_3;
assign _7 = ~(_2 | _15);
assign _14 = ~_5;
assign _8 = ~(_1 | _16);
assign _17 = ~_7;
assign _6 = ~(_13 | _14);
assign _18 = ~_8;
assign _9 = ~(_7 | _8);
assign _10 = ~(_17 | _18);
assign _11 = ~(_9 | _10);
assign _12 = ~(_6 | _11);
assign _4 = _12;
endmodule
