module gate(_0, _1, _2, _3, _594);
input _0, _1, _2, _3;
output _594;
wire _582, _583, _584, _585, _586, _587, _588, _589, _590, _591, _592, _593;
assign _584 = ~_0;
assign _583 = ~_1;
assign _586 = ~(_0 | _1);
assign _582 = ~_3;
assign _590 = ~(_2 | _584);
assign _587 = ~_586;
assign _585 = ~(_2 | _582);
assign _589 = ~(_582 | _583);
assign _588 = ~(_585 | _587);
assign _591 = ~(_589 | _590);
assign _592 = ~_591;
assign _593 = ~(_588 | _592);
assign _594 = _593;
endmodule
