module gate(_0, _1, _2, _3, _1299);
input _0, _1, _2, _3;
output _1299;
wire _1289, _1290, _1291, _1292, _1293, _1294, _1295, _1296, _1297, _1298;
assign _1291 = ~(_0 | _1);
assign _1290 = ~_2;
assign _1289 = ~_3;
assign _1292 = ~(_1290 | _1291);
assign _1294 = ~(_0 | _1290);
assign _1293 = ~_1292;
assign _1295 = ~(_1 | _1294);
assign _1297 = ~(_1289 | _1293);
assign _1296 = ~(_3 | _1295);
assign _1298 = ~(_1296 | _1297);
assign _1299 = _1298;
endmodule
