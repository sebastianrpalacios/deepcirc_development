module gate(_0, _1, _2, _3, _1230);
input _0, _1, _2, _3;
output _1230;
wire _1214, _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226, _1227, _1228, _1229;
assign _1217 = ~_0;
assign _1216 = ~_1;
assign _1215 = ~_2;
assign _1225 = ~(_1 | _2);
assign _1214 = ~_3;
assign _1221 = ~(_3 | _1215);
assign _1218 = ~(_2 | _1214);
assign _1222 = ~(_1217 | _1221);
assign _1219 = ~(_1216 | _1218);
assign _1223 = ~_1222;
assign _1226 = ~(_1222 | _1225);
assign _1220 = ~_1219;
assign _1227 = ~_1226;
assign _1224 = ~(_1220 | _1223);
assign _1228 = ~(_1219 | _1227);
assign _1229 = ~(_1224 | _1228);
assign _1230 = _1229;
endmodule
