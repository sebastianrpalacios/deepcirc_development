module m0x33 (input in2, in1, in3, output out);



endmodule
