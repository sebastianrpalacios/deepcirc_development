module gate(_0, _1, _2, _3, _248);
input _0, _1, _2, _3;
output _248;
wire _230, _231, _232, _233, _234, _235, _236, _237, _238, _239, _240, _241, _242, _243, _244, _245, _246, _247;
assign _233 = ~_0;
assign _231 = ~_1;
assign _232 = ~_2;
assign _230 = ~_3;
assign _236 = ~(_2 | _233);
assign _234 = ~(_3 | _231);
assign _241 = ~(_0 | _232);
assign _239 = ~(_1 | _230);
assign _237 = ~_236;
assign _235 = ~_234;
assign _244 = ~(_234 | _236);
assign _242 = ~_241;
assign _240 = ~_239;
assign _238 = ~(_235 | _237);
assign _245 = ~_244;
assign _243 = ~(_240 | _242);
assign _246 = ~(_243 | _245);
assign _247 = ~(_238 | _246);
assign _248 = _247;
endmodule
