module gate(_0, _1, _2, _3, _1119);
input _0, _1, _2, _3;
output _1119;
wire _1106, _1107, _1108, _1109, _1110, _1111, _1112, _1113, _1114, _1115, _1116;
assign _1109 = ~_0;
assign _1107 = ~_1;
assign _1108 = ~_2;
assign _1106 = ~_3;
assign _1113 = ~(_2 | _1109);
assign _1110 = ~(_0 | _1108);
assign _1111 = ~(_1106 | _1110);
assign _1114 = ~(_1107 | _1110);
assign _1112 = ~(_1 | _1111);
assign _1115 = ~_1114;
assign _1116 = ~(_1113 | _1115);
assign _1119 = _1112 | _1116;
endmodule
