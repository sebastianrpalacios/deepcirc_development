module gate(_0, _1, _2, _3, _607);
input _0, _1, _2, _3;
output _607;
wire _595, _596, _597, _598, _599, _600, _601, _602, _603, _604, _605, _606;
assign _598 = ~_0;
assign _596 = ~_1;
assign _597 = ~_2;
assign _595 = ~_3;
assign _600 = ~(_597 | _598);
assign _599 = ~(_2 | _595);
assign _601 = ~(_0 | _599);
assign _603 = ~(_599 | _600);
assign _602 = ~_601;
assign _604 = ~(_596 | _603);
assign _605 = ~(_1 | _602);
assign _606 = ~(_604 | _605);
assign _607 = _606;
endmodule
