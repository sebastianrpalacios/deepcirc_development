module m0x05 (input in2, in1, in3, output out);

	wire \$n6_0;
	wire \$n5_0;

	not (\$n5_0, in3);
	not (\$n6_0, in1);
	nor (out, \$n6_0, \$n5_0);

endmodule
