module gate(_0, _1, _2, _3, _1447);
input _0, _1, _2, _3;
output _1447;
wire _1433, _1434, _1435, _1436, _1437, _1438, _1439, _1440, _1441, _1442, _1443, _1444;
assign _1436 = ~_0;
assign _1435 = ~_1;
assign _1434 = ~_2;
assign _1433 = ~_3;
assign _1437 = ~(_3 | _1435);
assign _1440 = ~(_1434 | _1435);
assign _1442 = ~(_1 | _1433);
assign _1438 = ~(_1436 | _1437);
assign _1443 = ~(_2 | _1442);
assign _1439 = ~_1438;
assign _1441 = ~(_1438 | _1440);
assign _1444 = ~(_1439 | _1443);
assign _1447 = _1441 | _1444;
endmodule
