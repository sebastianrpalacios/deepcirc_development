module m0xAA (input in2, in1, in3, output out);


	not (out, in3);

endmodule
