module gate(_0, _1, _2, _3, _897);
input _0, _1, _2, _3;
output _897;
wire _884, _885, _886, _887, _888, _889, _890, _891, _892, _893, _894, _895, _896;
assign _887 = ~_0;
assign _885 = ~_1;
assign _886 = ~_2;
assign _884 = ~_3;
assign _888 = ~(_0 | _3);
assign _890 = ~(_884 | _887);
assign _889 = ~_888;
assign _893 = ~(_885 | _888);
assign _891 = ~(_888 | _890);
assign _894 = ~(_1 | _889);
assign _892 = ~(_886 | _891);
assign _895 = ~(_893 | _894);
assign _896 = ~(_892 | _895);
assign _897 = _896;
endmodule
