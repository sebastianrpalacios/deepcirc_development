module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _19, _20, _5, _6, _7, _8, _9;
assign _15 = ~_0;
assign _18 = ~_1;
assign _5 = ~(_0 | _1);
assign _17 = ~_2;
assign _16 = ~_3;
assign _14 = ~_5;
assign _11 = ~(_2 | _5);
assign _7 = ~(_15 | _16);
assign _6 = ~(_3 | _14);
assign _20 = ~_11;
assign _19 = ~_7;
assign _8 = ~(_6 | _7);
assign _10 = ~(_18 | _19);
assign _9 = ~(_8 | _17);
assign _12 = ~(_10 | _20);
assign _13 = ~(_9 | _12);
assign _4 = _13;
endmodule
