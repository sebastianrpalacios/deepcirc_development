module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _14, _15, _16, _17, _18, _19, _20, _21, _5, _6, _7, _8, _9;
assign _14 = ~_0;
assign _18 = ~_1;
assign _15 = ~_2;
assign _10 = ~(_1 | _2);
assign _16 = ~_3;
assign _5 = ~(_0 | _3);
assign _6 = ~(_14 | _15);
assign _21 = ~_10;
assign _20 = ~_5;
assign _8 = ~(_5 | _18);
assign _17 = ~_6;
assign _11 = ~(_20 | _21);
assign _19 = ~_8;
assign _7 = ~(_16 | _17);
assign _9 = ~(_7 | _19);
assign _4 = _9 | _11;
endmodule
