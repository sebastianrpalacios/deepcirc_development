module gate(_0, _1, _2, _3, _127);
input _0, _1, _2, _3;
output _127;
wire _118, _119, _120, _121, _122, _123, _124, _125, _126;
assign _118 = ~_1;
assign _119 = ~_2;
assign _122 = ~(_0 | _3);
assign _120 = ~(_3 | _118);
assign _123 = ~(_118 | _119);
assign _121 = ~(_2 | _120);
assign _124 = ~(_122 | _123);
assign _125 = ~_124;
assign _126 = ~(_121 | _125);
assign _127 = _126;
endmodule
