module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _15, _16, _17, _18, _19, _20, _21, _22, _23, _5, _6, _7, _8, _9;
assign _15 = ~_0;
assign _22 = ~_0;
assign _16 = ~_1;
assign _20 = ~_1;
assign _18 = ~_2;
assign _17 = ~_3;
assign _19 = ~_3;
assign _21 = ~_3;
assign _5 = ~(_15 | _16);
assign _8 = ~(_2 | _19);
assign _10 = ~(_20 | _21);
assign _6 = ~(_5 | _17);
assign _9 = ~(_1 | _8);
assign _11 = ~(_10 | _22);
assign _7 = ~(_6 | _18);
assign _23 = ~_11;
assign _12 = ~(_9 | _23);
assign _4 = _7 | _12;
endmodule
