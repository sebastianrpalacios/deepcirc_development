module gate(_0, _1, _2, _3, _283);
input _0, _1, _2, _3;
output _283;
wire _269, _270, _271, _272, _273, _274, _275, _276, _277, _278, _279, _280;
assign _272 = ~_0;
assign _271 = ~_1;
assign _270 = ~_2;
assign _269 = ~_3;
assign _278 = ~(_2 | _272);
assign _273 = ~(_269 | _270);
assign _276 = ~(_269 | _272);
assign _274 = ~_273;
assign _277 = ~(_271 | _276);
assign _275 = ~(_1 | _274);
assign _279 = ~(_277 | _278);
assign _280 = ~_279;
assign _283 = _275 | _280;
endmodule
