module gate(_0, _1, _2, _3, _1345);
input _0, _1, _2, _3;
output _1345;
wire _1333, _1334, _1335, _1336, _1337, _1338, _1339, _1340, _1341, _1342, _1343, _1344;
assign _1334 = ~_1;
assign _1335 = ~_2;
assign _1333 = ~_3;
assign _1337 = ~(_3 | _1334);
assign _1336 = ~(_0 | _1335);
assign _1341 = ~(_1333 | _1335);
assign _1338 = ~_1337;
assign _1339 = ~(_1334 | _1336);
assign _1342 = ~(_0 | _1341);
assign _1340 = ~(_1336 | _1338);
assign _1343 = ~(_1339 | _1342);
assign _1344 = ~(_1340 | _1343);
assign _1345 = _1344;
endmodule
