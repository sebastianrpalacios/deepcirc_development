module gate(_0, _1, _2, _3, _1176);
input _0, _1, _2, _3;
output _1176;
wire _1164, _1165, _1166, _1167, _1168, _1169, _1170, _1171, _1172, _1173, _1174, _1175;
assign _1166 = ~_0;
assign _1164 = ~_1;
assign _1165 = ~_2;
assign _1167 = ~(_0 | _2);
assign _1170 = ~(_1 | _2);
assign _1172 = ~(_1165 | _1166);
assign _1168 = ~(_3 | _1167);
assign _1173 = ~(_1164 | _1172);
assign _1169 = ~_1168;
assign _1171 = ~(_1168 | _1170);
assign _1174 = ~(_1169 | _1173);
assign _1175 = ~(_1171 | _1174);
assign _1176 = _1175;
endmodule
