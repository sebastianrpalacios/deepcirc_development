module gate(_0, _1, _2, _3, _761);
input _0, _1, _2, _3;
output _761;
wire _747, _748, _749, _750, _751, _752, _753, _754, _755, _756, _757, _758, _759, _760;
assign _748 = ~_1;
assign _749 = ~_2;
assign _747 = ~_3;
assign _753 = ~(_2 | _3);
assign _750 = ~(_1 | _749);
assign _752 = ~(_748 | _749);
assign _751 = ~(_2 | _747);
assign _756 = ~(_747 | _749);
assign _755 = ~(_752 | _753);
assign _754 = ~(_750 | _751);
assign _757 = ~(_0 | _756);
assign _759 = ~(_0 | _755);
assign _758 = ~(_754 | _757);
assign _760 = ~(_758 | _759);
assign _761 = _760;
endmodule
