module m0x55 (input in2, in1, in3, output out);



endmodule
