module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _19, _20, _5, _6, _7, _8, _9;
assign _15 = ~_0;
assign _13 = ~_1;
assign _17 = ~_1;
assign _14 = ~_2;
assign _5 = ~(_1 | _2);
assign _18 = ~_3;
assign _7 = ~(_3 | _15);
assign _9 = ~(_0 | _17);
assign _6 = ~(_13 | _14);
assign _16 = ~_7;
assign _19 = ~_9;
assign _8 = ~(_6 | _16);
assign _10 = ~(_18 | _19);
assign _11 = ~(_5 | _8);
assign _20 = ~_11;
assign _12 = ~(_10 | _20);
assign _4 = _12;
endmodule
