module gate(_0, _1, _2, _3, _527);
input _0, _1, _2, _3;
output _527;
wire _515, _516, _517, _518, _519, _520, _521, _522, _523, _524, _525, _526;
assign _518 = ~_0;
assign _516 = ~_1;
assign _517 = ~_2;
assign _515 = ~_3;
assign _519 = ~(_2 | _516);
assign _520 = ~(_1 | _517);
assign _521 = ~(_515 | _520);
assign _522 = ~_521;
assign _523 = ~(_518 | _521);
assign _524 = ~(_0 | _522);
assign _525 = ~(_523 | _524);
assign _526 = ~(_519 | _525);
assign _527 = _526;
endmodule
