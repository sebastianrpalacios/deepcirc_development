module gate(_0, _1, _2, _3, _620);
input _0, _1, _2, _3;
output _620;
wire _608, _609, _610, _611, _612, _613, _614, _615, _616, _617, _618, _619;
assign _610 = ~_0;
assign _609 = ~_1;
assign _608 = ~_3;
assign _613 = ~(_1 | _610);
assign _611 = ~(_0 | _609);
assign _612 = ~_611;
assign _614 = ~(_611 | _613);
assign _616 = ~(_608 | _611);
assign _617 = ~(_3 | _612);
assign _615 = ~(_2 | _614);
assign _618 = ~(_616 | _617);
assign _619 = ~(_615 | _618);
assign _620 = _619;
endmodule
