module gate(_0, _1, _2, _3, _1201);
input _0, _1, _2, _3;
output _1201;
wire _1190, _1191, _1192, _1193, _1194, _1195, _1196, _1197, _1198, _1199, _1200;
assign _1192 = ~_0;
assign _1193 = ~(_0 | _1);
assign _1191 = ~_2;
assign _1190 = ~_3;
assign _1194 = ~(_3 | _1193);
assign _1196 = ~(_1190 | _1192);
assign _1195 = ~_1194;
assign _1197 = ~(_1193 | _1196);
assign _1199 = ~(_2 | _1195);
assign _1198 = ~(_1191 | _1197);
assign _1200 = ~(_1198 | _1199);
assign _1201 = _1200;
endmodule
