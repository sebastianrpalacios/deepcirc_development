module gate(_0, _1, _2, _3, _1028);
input _0, _1, _2, _3;
output _1028;
wire _1012, _1013, _1014, _1015, _1016, _1017, _1018, _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027;
assign _1015 = ~_0;
assign _1014 = ~_1;
assign _1013 = ~_2;
assign _1012 = ~_3;
assign _1016 = ~(_1 | _1015);
assign _1021 = ~(_2 | _1014);
assign _1018 = ~(_3 | _1013);
assign _1017 = ~_1016;
assign _1024 = ~(_1012 | _1016);
assign _1022 = ~_1021;
assign _1019 = ~_1018;
assign _1023 = ~(_0 | _1022);
assign _1020 = ~(_1017 | _1019);
assign _1025 = ~(_1020 | _1024);
assign _1026 = ~_1025;
assign _1027 = ~(_1023 | _1026);
assign _1028 = _1027;
endmodule
