module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _16, _17, _18, _19, _20, _21, _5, _6, _7, _8, _9;
assign _18 = ~_0;
assign _19 = ~_1;
assign _16 = ~_2;
assign _9 = ~(_0 | _2);
assign _17 = ~_3;
assign _20 = ~_3;
assign _5 = ~(_2 | _3);
assign _10 = ~(_1 | _9);
assign _6 = ~(_16 | _17);
assign _11 = ~(_19 | _20);
assign _7 = ~(_5 | _6);
assign _12 = ~(_5 | _11);
assign _8 = ~(_7 | _18);
assign _21 = ~_12;
assign _13 = ~(_10 | _21);
assign _4 = _8 | _13;
endmodule
