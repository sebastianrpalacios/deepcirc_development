module gate(_0, _1, _2, _3, _339);
input _0, _1, _2, _3;
output _339;
wire _329, _330, _331, _332, _333, _334, _335, _336, _337, _338;
assign _331 = ~_0;
assign _329 = ~_1;
assign _330 = ~_2;
assign _335 = ~(_1 | _2);
assign _332 = ~(_330 | _331);
assign _336 = ~(_3 | _335);
assign _333 = ~_332;
assign _337 = ~(_332 | _336);
assign _334 = ~(_329 | _333);
assign _338 = ~(_334 | _337);
assign _339 = _338;
endmodule
