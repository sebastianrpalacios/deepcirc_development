module gate(_0, _1, _2, _3, _141);
input _0, _1, _2, _3;
output _141;
wire _128, _129, _130, _131, _132, _133, _134, _135, _136, _137, _138, _139, _140;
assign _130 = ~_0;
assign _128 = ~_1;
assign _129 = ~_2;
assign _134 = ~(_0 | _2);
assign _131 = ~(_2 | _3);
assign _135 = ~(_1 | _3);
assign _133 = ~(_129 | _130);
assign _132 = ~(_128 | _131);
assign _136 = ~(_134 | _135);
assign _137 = ~_136;
assign _138 = ~(_133 | _137);
assign _139 = ~_138;
assign _140 = ~(_132 | _139);
assign _141 = _140;
endmodule
