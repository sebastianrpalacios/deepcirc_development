module gate(_0, _1, _2, _3, _410);
input _0, _1, _2, _3;
output _410;
wire _396, _397, _398, _399, _400, _401, _402, _403, _404, _405, _406, _407;
assign _399 = ~_0;
assign _397 = ~_1;
assign _398 = ~_2;
assign _396 = ~_3;
assign _404 = ~(_2 | _397);
assign _400 = ~(_1 | _398);
assign _401 = ~(_396 | _397);
assign _405 = ~(_399 | _400);
assign _402 = ~(_400 | _401);
assign _406 = ~_405;
assign _403 = ~(_0 | _402);
assign _407 = ~(_404 | _406);
assign _410 = _403 | _407;
endmodule
