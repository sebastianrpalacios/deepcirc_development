module gate(_0, _1, _2, _3, _1213);
input _0, _1, _2, _3;
output _1213;
wire _1202, _1203, _1204, _1205, _1206, _1207, _1208, _1209, _1210, _1211, _1212;
assign _1205 = ~_0;
assign _1203 = ~_1;
assign _1204 = ~_2;
assign _1202 = ~_3;
assign _1206 = ~(_0 | _3);
assign _1207 = ~(_2 | _1203);
assign _1208 = ~(_1 | _1204);
assign _1209 = ~(_1202 | _1205);
assign _1210 = ~(_1207 | _1209);
assign _1211 = ~(_1206 | _1210);
assign _1212 = ~(_1208 | _1211);
assign _1213 = _1212;
endmodule
