module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _5, _6, _7, _8, _9;
assign _18 = ~_0;
assign _14 = ~_1;
assign _15 = ~_2;
assign _17 = ~_3;
assign _10 = ~(_1 | _18);
assign _5 = ~(_0 | _14);
assign _9 = ~(_1 | _17);
assign _11 = ~(_3 | _10);
assign _16 = ~_5;
assign _6 = ~(_5 | _15);
assign _12 = ~(_9 | _11);
assign _7 = ~(_2 | _16);
assign _8 = ~(_6 | _7);
assign _13 = ~(_8 | _12);
assign _4 = _13;
endmodule
