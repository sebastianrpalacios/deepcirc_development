module gate(_0, _1, _2, _3, _633);
input _0, _1, _2, _3;
output _633;
wire _621, _622, _623, _624, _625, _626, _627, _628, _629, _630, _631, _632;
assign _624 = ~_0;
assign _622 = ~_1;
assign _623 = ~_2;
assign _621 = ~_3;
assign _628 = ~(_622 | _623);
assign _625 = ~(_1 | _621);
assign _626 = ~_625;
assign _629 = ~(_0 | _625);
assign _627 = ~(_624 | _626);
assign _630 = ~_629;
assign _631 = ~(_628 | _630);
assign _632 = ~(_627 | _631);
assign _633 = _632;
endmodule
