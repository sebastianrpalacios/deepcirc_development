module gate(_0, _1, _2, _3, _703);
input _0, _1, _2, _3;
output _703;
wire _691, _692, _693, _694, _695, _696, _697, _698, _699, _700, _701, _702;
assign _694 = ~_0;
assign _692 = ~_1;
assign _698 = ~(_0 | _1);
assign _693 = ~_2;
assign _691 = ~_3;
assign _695 = ~(_692 | _693);
assign _696 = ~(_694 | _695);
assign _699 = ~(_695 | _698);
assign _697 = ~_696;
assign _700 = ~(_3 | _699);
assign _701 = ~(_691 | _697);
assign _702 = ~(_700 | _701);
assign _703 = _702;
endmodule
