module gate(_0, _1, _2, _3, _351);
input _0, _1, _2, _3;
output _351;
wire _340, _341, _342, _343, _344, _345, _346, _347, _348, _349, _350;
assign _342 = ~_0;
assign _341 = ~_1;
assign _340 = ~_2;
assign _346 = ~(_1 | _2);
assign _343 = ~(_340 | _341);
assign _347 = ~(_3 | _346);
assign _344 = ~(_342 | _343);
assign _345 = ~_344;
assign _348 = ~(_344 | _347);
assign _349 = ~(_3 | _345);
assign _350 = ~(_348 | _349);
assign _351 = _350;
endmodule
