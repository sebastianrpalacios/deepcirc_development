module gate(_0, _1, _2, _3, _1189);
input _0, _1, _2, _3;
output _1189;
wire _1177, _1178, _1179, _1180, _1181, _1182, _1183, _1184, _1185, _1186, _1187, _1188;
assign _1179 = ~_0;
assign _1178 = ~_1;
assign _1180 = ~_2;
assign _1177 = ~_3;
assign _1183 = ~(_3 | _1178);
assign _1181 = ~(_1177 | _1178);
assign _1182 = ~(_1177 | _1179);
assign _1186 = ~(_1179 | _1181);
assign _1184 = ~(_1182 | _1183);
assign _1187 = ~(_1180 | _1186);
assign _1185 = ~(_2 | _1184);
assign _1188 = ~(_1185 | _1187);
assign _1189 = _1188;
endmodule
