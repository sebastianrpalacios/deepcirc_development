module gate(_0, _1, _2, _3, _567);
input _0, _1, _2, _3;
output _567;
wire _556, _557, _558, _559, _560, _561, _562, _563, _564;
assign _558 = ~_0;
assign _557 = ~_1;
assign _556 = ~_2;
assign _559 = ~(_556 | _557);
assign _561 = ~(_0 | _556);
assign _563 = ~(_1 | _556);
assign _560 = ~(_558 | _559);
assign _562 = ~(_3 | _561);
assign _564 = ~(_562 | _563);
assign _567 = _560 | _564;
endmodule
