module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _17, _18, _5, _6, _7, _8, _9;
assign _13 = ~_0;
assign _16 = ~_1;
assign _14 = ~_3;
assign _5 = ~(_3 | _13);
assign _6 = ~(_0 | _14);
assign _15 = ~_5;
assign _7 = ~(_5 | _6);
assign _8 = ~(_2 | _15);
assign _18 = ~_7;
assign _9 = ~(_7 | _16);
assign _11 = ~(_1 | _18);
assign _17 = ~_9;
assign _10 = ~(_8 | _17);
assign _12 = ~(_10 | _11);
assign _4 = _12;
endmodule
