module gate(_0, _1, _2, _3, _1045);
input _0, _1, _2, _3;
output _1045;
wire _1029, _1030, _1031, _1032, _1033, _1034, _1035, _1036, _1037, _1038, _1039, _1040, _1041, _1042;
assign _1032 = ~_0;
assign _1031 = ~_1;
assign _1030 = ~_2;
assign _1029 = ~_3;
assign _1036 = ~(_2 | _1031);
assign _1033 = ~(_1 | _1030);
assign _1038 = ~(_1029 | _1031);
assign _1037 = ~(_3 | _1036);
assign _1034 = ~_1033;
assign _1039 = ~_1038;
assign _1035 = ~(_1032 | _1034);
assign _1040 = ~(_0 | _1039);
assign _1041 = ~(_1037 | _1040);
assign _1042 = ~_1041;
assign _1045 = _1035 | _1042;
endmodule
