module m0x88 (input in2, in1, in3, output out);


	nor (out, in2, in3);

endmodule
