module gate(_0, _1, _2, _3, _674);
input _0, _1, _2, _3;
output _674;
wire _660, _661, _662, _663, _664, _665, _666, _667, _668, _669, _670, _671;
assign _661 = ~_0;
assign _660 = ~_1;
assign _662 = ~(_0 | _1);
assign _665 = ~(_1 | _661);
assign _669 = ~(_2 | _661);
assign _663 = ~(_660 | _661);
assign _664 = ~(_0 | _660);
assign _670 = ~(_3 | _669);
assign _666 = ~(_662 | _663);
assign _667 = ~(_664 | _665);
assign _671 = ~(_666 | _670);
assign _668 = ~(_3 | _667);
assign _674 = _668 | _671;
endmodule
