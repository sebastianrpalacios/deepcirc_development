module gate(_0, _1, _2, _3, _802);
input _0, _1, _2, _3;
output _802;
wire _788, _789, _790, _791, _792, _793, _794, _795, _796, _797, _798, _799, _800, _801;
assign _789 = ~_0;
assign _788 = ~_1;
assign _790 = ~_2;
assign _794 = ~(_1 | _2);
assign _795 = ~(_788 | _789);
assign _791 = ~(_788 | _790);
assign _799 = ~(_0 | _794);
assign _796 = ~(_794 | _795);
assign _792 = ~(_3 | _791);
assign _797 = ~_796;
assign _793 = ~_792;
assign _798 = ~(_792 | _797);
assign _800 = ~(_793 | _799);
assign _801 = ~(_798 | _800);
assign _802 = _801;
endmodule
