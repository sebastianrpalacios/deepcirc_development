module gate(_0, _1, _2, _3, _1407);
input _0, _1, _2, _3;
output _1407;
wire _1396, _1397, _1398, _1399, _1400, _1401, _1402, _1403, _1404, _1405, _1406;
assign _1398 = ~_0;
assign _1397 = ~_1;
assign _1403 = ~(_1 | _2);
assign _1396 = ~_3;
assign _1400 = ~(_0 | _1397);
assign _1404 = ~_1403;
assign _1399 = ~(_2 | _1396);
assign _1401 = ~_1400;
assign _1405 = ~(_1398 | _1404);
assign _1402 = ~(_1399 | _1401);
assign _1406 = ~(_1402 | _1405);
assign _1407 = _1406;
endmodule
