module gate(_0, _1, _2, _3, _297);
input _0, _1, _2, _3;
output _297;
wire _284, _285, _286, _287, _288, _289, _290, _291, _292, _293, _294;
assign _286 = ~_0;
assign _285 = ~_1;
assign _287 = ~_2;
assign _284 = ~_3;
assign _288 = ~(_3 | _287);
assign _289 = ~(_2 | _284);
assign _290 = ~_289;
assign _292 = ~(_285 | _289);
assign _291 = ~(_1 | _290);
assign _293 = ~(_291 | _292);
assign _294 = ~(_286 | _293);
assign _297 = _288 | _294;
endmodule
