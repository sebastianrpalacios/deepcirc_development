module gate(_0, _1, _2, _3, _204);
input _0, _1, _2, _3;
output _204;
wire _192, _193, _194, _195, _196, _197, _198, _199, _200, _201;
assign _193 = ~_1;
assign _194 = ~_2;
assign _198 = ~(_1 | _2);
assign _192 = ~_3;
assign _195 = ~(_193 | _194);
assign _196 = ~_195;
assign _199 = ~(_195 | _198);
assign _197 = ~(_0 | _196);
assign _200 = ~_199;
assign _201 = ~(_192 | _200);
assign _204 = _197 | _201;
endmodule
