module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _14, _15, _16, _17, _18, _19, _5, _6, _7, _8, _9;
assign _15 = ~_0;
assign _14 = ~_1;
assign _17 = ~_2;
assign _16 = ~_3;
assign _5 = ~(_3 | _14);
assign _7 = ~(_1 | _16);
assign _6 = ~(_5 | _15);
assign _8 = ~(_5 | _7);
assign _18 = ~_8;
assign _9 = ~(_8 | _17);
assign _10 = ~(_2 | _18);
assign _11 = ~(_6 | _9);
assign _19 = ~_11;
assign _4 = _10 | _19;
endmodule
