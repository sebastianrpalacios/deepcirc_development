module gate(_0, _1, _2, _3, _690);
input _0, _1, _2, _3;
output _690;
wire _675, _676, _677, _678, _679, _680, _681, _682, _683, _684, _685, _686, _687, _688, _689;
assign _677 = ~_0;
assign _676 = ~_1;
assign _678 = ~_2;
assign _675 = ~_3;
assign _682 = ~(_1 | _3);
assign _685 = ~(_1 | _678);
assign _679 = ~(_675 | _676);
assign _683 = ~_682;
assign _686 = ~(_677 | _685);
assign _680 = ~_679;
assign _684 = ~(_0 | _683);
assign _681 = ~(_2 | _680);
assign _687 = ~(_684 | _686);
assign _688 = ~_687;
assign _689 = ~(_681 | _688);
assign _690 = _689;
endmodule
