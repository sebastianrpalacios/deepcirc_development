module gate(_0, _1, _2, _3, _1105);
input _0, _1, _2, _3;
output _1105;
wire _1088, _1089, _1090, _1091, _1092, _1093, _1094, _1095, _1096, _1097, _1098, _1099, _1100, _1101, _1102;
assign _1091 = ~_0;
assign _1089 = ~_1;
assign _1090 = ~_2;
assign _1097 = ~(_1 | _2);
assign _1088 = ~_3;
assign _1092 = ~(_3 | _1091);
assign _1094 = ~(_1089 | _1090);
assign _1098 = ~_1097;
assign _1093 = ~_1092;
assign _1095 = ~_1094;
assign _1100 = ~(_1092 | _1094);
assign _1099 = ~(_1088 | _1098);
assign _1096 = ~(_1093 | _1095);
assign _1101 = ~_1100;
assign _1102 = ~(_1099 | _1101);
assign _1105 = _1096 | _1102;
endmodule
