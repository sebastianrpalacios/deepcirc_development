module gate(_0, _1, _2, _3, _774);
input _0, _1, _2, _3;
output _774;
wire _762, _763, _764, _765, _766, _767, _768, _769, _770, _771, _772, _773;
assign _764 = ~_1;
assign _763 = ~_2;
assign _762 = ~_3;
assign _767 = ~(_0 | _764);
assign _765 = ~(_0 | _763);
assign _768 = ~(_762 | _767);
assign _771 = ~(_763 | _767);
assign _766 = ~(_1 | _765);
assign _769 = ~_768;
assign _772 = ~(_3 | _771);
assign _770 = ~(_766 | _769);
assign _773 = ~(_770 | _772);
assign _774 = _773;
endmodule
