module m0x4C (input in2, in1, in3, output out);

	wire \$new_n5__0;

	nor (\$new_n5__0, in1, in3);
	nor (out, \$new_n5__0, in2);

endmodule
