module gate(_0, _1, _2, _3, _541);
input _0, _1, _2, _3;
output _541;
wire _528, _529, _530, _531, _532, _533, _534, _535, _536, _537, _538, _539, _540;
assign _530 = ~_0;
assign _529 = ~_1;
assign _531 = ~_2;
assign _528 = ~_3;
assign _536 = ~(_1 | _3);
assign _533 = ~(_2 | _530);
assign _537 = ~(_2 | _529);
assign _532 = ~(_0 | _531);
assign _538 = ~(_536 | _537);
assign _534 = ~(_532 | _533);
assign _539 = ~(_533 | _538);
assign _535 = ~(_528 | _534);
assign _540 = ~(_535 | _539);
assign _541 = _540;
endmodule
