module gate(_0, _1, _2, _3, _1432);
input _0, _1, _2, _3;
output _1432;
wire _1423, _1424, _1425, _1426, _1427, _1428, _1429, _1430, _1431;
assign _1425 = ~_0;
assign _1424 = ~_1;
assign _1423 = ~_3;
assign _1426 = ~(_2 | _1424);
assign _1430 = ~(_3 | _1424);
assign _1427 = ~(_1423 | _1425);
assign _1428 = ~_1427;
assign _1429 = ~(_1426 | _1428);
assign _1431 = ~(_1429 | _1430);
assign _1432 = _1431;
endmodule
