module gate(_0, _1, _2, _3, _328);
input _0, _1, _2, _3;
output _328;
wire _316, _317, _318, _319, _320, _321, _322, _323, _324, _325, _326, _327;
assign _317 = ~_1;
assign _318 = ~_2;
assign _316 = ~_3;
assign _323 = ~(_0 | _317);
assign _319 = ~(_3 | _318);
assign _322 = ~(_2 | _316);
assign _324 = ~_323;
assign _320 = ~_319;
assign _325 = ~(_322 | _324);
assign _321 = ~(_0 | _320);
assign _326 = ~(_1 | _321);
assign _327 = ~(_325 | _326);
assign _328 = _327;
endmodule
