module m0xA0 (input in2, in1, in3, output out);


	nor (out, in1, in3);

endmodule
