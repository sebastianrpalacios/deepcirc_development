module gate(_0, _1, _2, _3, _932);
input _0, _1, _2, _3;
output _932;
wire _920, _921, _922, _923, _924, _925, _926, _927, _928, _929, _930, _931;
assign _923 = ~_0;
assign _921 = ~_1;
assign _922 = ~_2;
assign _924 = ~(_1 | _2);
assign _920 = ~_3;
assign _925 = ~(_921 | _923);
assign _928 = ~(_0 | _922);
assign _926 = ~(_924 | _925);
assign _929 = ~(_920 | _928);
assign _927 = ~_926;
assign _930 = ~(_3 | _927);
assign _931 = ~(_929 | _930);
assign _932 = _931;
endmodule
