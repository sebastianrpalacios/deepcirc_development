module gate(_0, _1, _2, _3, _171);
input _0, _1, _2, _3;
output _171;
wire _156, _157, _158, _159, _160, _161, _162, _163, _164, _165, _166, _167, _168, _169, _170;
assign _159 = ~_0;
assign _157 = ~_1;
assign _158 = ~_2;
assign _156 = ~_3;
assign _163 = ~(_1 | _3);
assign _166 = ~(_2 | _159);
assign _161 = ~(_3 | _157);
assign _167 = ~(_0 | _158);
assign _160 = ~(_1 | _156);
assign _162 = ~(_156 | _157);
assign _164 = ~(_160 | _161);
assign _165 = ~(_162 | _163);
assign _169 = ~(_164 | _167);
assign _168 = ~(_165 | _166);
assign _170 = ~(_168 | _169);
assign _171 = _170;
endmodule
