module gate(_0, _1, _2, _3, _4);
input _0, _1, _2, _3;
output _4;
wire _10, _11, _12, _13, _14, _15, _16, _19, _20, _21, _22, _23, _24, _25, _26, _5, _6, _7, _8, _9;
assign _19 = ~_0;
assign _23 = ~_1;
assign _8 = ~(_0 | _1);
assign _21 = ~_2;
assign _24 = ~_2;
assign _20 = ~_3;
assign _5 = ~(_1 | _19);
assign _13 = ~(_0 | _23);
assign _22 = ~_8;
assign _9 = ~(_8 | _21);
assign _6 = ~(_0 | _20);
assign _15 = ~(_3 | _5);
assign _25 = ~_13;
assign _10 = ~(_2 | _22);
assign _7 = ~(_5 | _6);
assign _26 = ~_15;
assign _14 = ~(_24 | _25);
assign _11 = ~(_9 | _10);
assign _16 = ~(_14 | _26);
assign _12 = ~(_7 | _11);
assign _4 = _12 | _16;
endmodule
