module gate(_0, _1, _2, _3, _452);
input _0, _1, _2, _3;
output _452;
wire _437, _438, _439, _440, _441, _442, _443, _444, _445, _446, _447, _448, _449, _450, _451;
assign _440 = ~_0;
assign _438 = ~_1;
assign _439 = ~_2;
assign _443 = ~(_1 | _2);
assign _437 = ~_3;
assign _441 = ~(_3 | _440);
assign _444 = ~(_438 | _439);
assign _446 = ~(_437 | _438);
assign _442 = ~_441;
assign _447 = ~_446;
assign _445 = ~(_442 | _444);
assign _448 = ~(_0 | _447);
assign _449 = ~(_445 | _448);
assign _450 = ~_449;
assign _451 = ~(_443 | _450);
assign _452 = _451;
endmodule
