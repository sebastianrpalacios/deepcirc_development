module gate(_0, _1, _2, _3, _502);
input _0, _1, _2, _3;
output _502;
wire _486, _487, _488, _489, _490, _491, _492, _493, _494, _495, _496, _497, _498, _499;
assign _488 = ~_0;
assign _497 = ~(_0 | _1);
assign _487 = ~_2;
assign _486 = ~_3;
assign _489 = ~(_1 | _3);
assign _498 = ~_497;
assign _492 = ~(_2 | _486);
assign _490 = ~_489;
assign _493 = ~_492;
assign _494 = ~(_488 | _492);
assign _491 = ~(_487 | _490);
assign _499 = ~(_493 | _498);
assign _495 = ~_494;
assign _496 = ~(_491 | _495);
assign _502 = _496 | _499;
endmodule
